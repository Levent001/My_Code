`timescale 1ns / 1ps
`include "./axi_stream_insert_header.v"
module test_module;

    parameter PERIOD = 10;
    parameter DATA_WD = 32;
    parameter DATA_BYTE_WD = DATA_WD / 8;
    parameter BYTE_CNT_WD = $clog2(DATA_BYTE_WD);
    parameter tb_datain_depth = 4;

    // axi_stream_insert_header Inputs
    reg                       clk = 1;
    reg                       rst_n = 0;
    reg                       valid_in = 0;
    reg  [     DATA_WD-1 : 0] data_in = 0;
    reg  [DATA_BYTE_WD-1 : 0] keep_in = 0;
    reg                       ready_out = 1;
    reg                       valid_insert = 0;
    reg  [     DATA_WD-1 : 0] header_insert = 0;
    reg  [DATA_BYTE_WD-1 : 0] keep_insert = 0;
    reg  [   BYTE_CNT_WD : 0] byte_insert_cnt = 0;

    // axi_stream_insert_header Outputs
    wire                      ready_in;
    wire                      valid_out;
    wire [     DATA_WD-1 : 0] data_out;
    wire [DATA_BYTE_WD-1 : 0] keep_out;
    wire                      last_out;
    wire                      ready_insert;
    reg                       last_in = 0;
    reg valid_insert_tmp;
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n)
            valid_insert_tmp <= 0;
        else begin
            valid_insert_tmp <= ready_in;
        end
    end

    initial begin
        forever #(PERIOD / 2) clk = ~clk;
    end

    initial begin
        #PERIOD
        rst_n = 1;

        #PERIOD 
        valid_insert = 1;
        ready_out = 1;
        header_insert = 32'hFFEEDDCC;
        keep_insert = 4'b0111;
        
        #PERIOD
        valid_insert = 0;
        valid_in = 1;
        data_in = 32'hAABBCCDD;
        keep_in = 4'b1111;
        #PERIOD
        data_in = 32'hEEFF0011;
        keep_in = 4'b1111;
        #PERIOD
        data_in = 32'h22334455;
        keep_in = 4'b1111;
        #PERIOD
        data_in = 32'h66778899;
        keep_in = 4'b1111;
        #PERIOD
        data_in = 32'hAABB0000;
        keep_in = 4'b1100;
        last_in = 1;
    end

    axi_stream_insert_header #(
        .DATA_WD     (DATA_WD),
        .DATA_BYTE_WD(DATA_BYTE_WD)
    ) u_axi_stream_insert_header (
        .clk         (clk),
        .rst_n       (rst_n),
        .valid_in    (valid_in),
        .data_in     (data_in[DATA_WD-1 : 0]),
        .keep_in     (keep_in[DATA_BYTE_WD-1 : 0]),
        .last_in     (last_in),
        .ready_out   (ready_out),
        .valid_insert(valid_insert),
        .header_insert (header_insert[DATA_WD-1 : 0]),
        .keep_insert (keep_insert[DATA_BYTE_WD-1 : 0]),

        .ready_in    (ready_in),
        .valid_out   (valid_out),
        .data_out    (data_out[DATA_WD-1 : 0]),
        .keep_out    (keep_out[DATA_BYTE_WD-1 : 0]),
        .last_out    (last_out),
        .ready_insert(ready_insert)
    );

    

////////////////////////////////////////////////////////////
    initial begin
        $dumpfile("wave.vcd");  //生成的vcd文件名称
        $dumpvars(0, test_module);  //tb模块名称
        #20000 $finish;
    end
////////////////////////////////////////////////////////////
endmodule
